CONFIG_TARGET:cfg_core_arm
CONFIG_IRQ2EN:0
CFG_DCACHE_LSZ:4
CFG_ICACHE_REPL:cfg_repl_rnd
CFG_DCACHE_ALLOCATE:0
CFG_DCACHE_ALGO:rnd
CFG_ICACHE_SZ:1
CFG_ICACHE_LOCK:0
CFG_ICACHE_LSZ:4
CFG_DCACHE_ASSO:1
CFG_DCACHE_TYPE:writethrough
CFG_DCACHE_LOCK:0
CFG_ICACHE_ASSO:1
CFG_DCACHE_REPL:cfg_repl_rnd
CFG_DCACHE_SZ:1
CFG_DCACHE_WB:2
CFG_ICACHE_ALGO:rnd
CONFIG_BOOT_SYSCLK:25000000
CONFIG_IRQ2EN:0
CONFIG_IRQ2CHAN:1
CONFIG_WDOG:0
